3
2 2 1 2 3 g  0x4de6f50  0x4de7fd0  0x4de7310 c  10 1 15 3 27 2
10 12 21 39 3 g  0x4de6420  0x4de64f0  0x4de65d0 c  7 1 34 2
12 6 3 11 3 g  0x4de6890  0x4de6bd0  0x4de6dd0  0x4de7410  0x4de7290  0x4de66d0  0x4de6910 c  2 3 14 3 6 3 2 3 2 3 14 3 14 3 6 3
1 1 10 2 0 g  0x4de8c50  0x4de9690  0x4de85d0  0x4de7510  0x4de9890  0x4de9990  0x4de9710 c  53 1 45 1 38 2
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
0
